-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Thu May 22 09:36:15 2014"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY sensordeled IS 
	PORT
	(
		Vaga1 :  IN  STD_LOGIC;
		Vaga2 :  IN  STD_LOGIC;
		Vaga3 :  IN  STD_LOGIC;
		Vaga4 :  IN  STD_LOGIC;
		Vaga5 :  IN  STD_LOGIC;
		Vaga6 :  IN  STD_LOGIC;
		Vaga7 :  IN  STD_LOGIC;
		Vaga8 :  IN  STD_LOGIC;
		Vaga9 :  IN  STD_LOGIC;
		Vaga11 :  IN  STD_LOGIC;
		Vaga10 :  IN  STD_LOGIC;
		Vaga12 :  IN  STD_LOGIC;
		Vaga13 :  IN  STD_LOGIC;
		Vaga14 :  IN  STD_LOGIC;
		Vaga15 :  IN  STD_LOGIC;
		Vaga16 :  IN  STD_LOGIC;
		Led_Vaga2 :  OUT  STD_LOGIC;
		Led_Vaga3 :  OUT  STD_LOGIC;
		Led_Vaga4 :  OUT  STD_LOGIC;
		Led_Vaga5 :  OUT  STD_LOGIC;
		Led_Vaga6 :  OUT  STD_LOGIC;
		Led_Vaga7 :  OUT  STD_LOGIC;
		Led_Vaga_Deficiente :  OUT  STD_LOGIC;
		Led_Vaga8 :  OUT  STD_LOGIC;
		Led_Vaga9 :  OUT  STD_LOGIC;
		Led_Vaga10 :  OUT  STD_LOGIC;
		Led_Vaga11 :  OUT  STD_LOGIC;
		Led_Vaga12 :  OUT  STD_LOGIC;
		Led_Vaga13 :  OUT  STD_LOGIC;
		Led_Vaga14 :  OUT  STD_LOGIC;
		Led_Vaga15 :  OUT  STD_LOGIC;
		pin_name1 :  OUT  STD_LOGIC;
		pin_name2 :  OUT  STD_LOGIC;
		pin_name3 :  OUT  STD_LOGIC;
		pin_name4 :  OUT  STD_LOGIC;
		Led_Vaga1 :  OUT  STD_LOGIC
	);
END sensordeled;

ARCHITECTURE bdf_type OF sensordeled IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \74283_0\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_0\: COMPONENT IS true;

COMPONENT \74283_1\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_1\: COMPONENT IS true;

COMPONENT \74283_10\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_10\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_10\: COMPONENT IS true;

COMPONENT \74283_11\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_11\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_11\: COMPONENT IS true;

COMPONENT \74283_12\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_12\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_12\: COMPONENT IS true;

COMPONENT \74283_13\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_13\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_13\: COMPONENT IS true;

COMPONENT \74283_2\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_2\: COMPONENT IS true;

COMPONENT \74283_3\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_3\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_3\: COMPONENT IS true;

COMPONENT \74283_4\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_4\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_4\: COMPONENT IS true;

COMPONENT \74283_5\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_5\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_5\: COMPONENT IS true;

COMPONENT \74283_6\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_6\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_6\: COMPONENT IS true;

COMPONENT \74283_7\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_7\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_7\: COMPONENT IS true;

COMPONENT \74283_8\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_8\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_8\: COMPONENT IS true;

COMPONENT \74283_9\
	PORT(CIN : IN STD_LOGIC;
		 A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 SUM4 : OUT STD_LOGIC;
		 SUM1 : OUT STD_LOGIC;
		 SUM2 : OUT STD_LOGIC;
		 SUM3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74283_9\: COMPONENT IS true;
ATTRIBUTE noopt OF \74283_9\: COMPONENT IS true;

SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;


BEGIN 
Led_Vaga2 <= Vaga2;
Led_Vaga3 <= Vaga3;
Led_Vaga4 <= Vaga4;
Led_Vaga5 <= Vaga5;
Led_Vaga6 <= Vaga6;
Led_Vaga7 <= Vaga7;
Led_Vaga_Deficiente <= Vaga16;
Led_Vaga8 <= Vaga8;
Led_Vaga9 <= Vaga9;
Led_Vaga10 <= Vaga10;
Led_Vaga11 <= Vaga11;
Led_Vaga12 <= Vaga12;
Led_Vaga13 <= Vaga13;
Led_Vaga14 <= Vaga14;
Led_Vaga15 <= Vaga15;
Led_Vaga1 <= Vaga1;
SYNTHESIZED_WIRE_7 <= '1';
SYNTHESIZED_WIRE_56 <= '1';
SYNTHESIZED_WIRE_113 <= '1';
SYNTHESIZED_WIRE_114 <= '1';
SYNTHESIZED_WIRE_115 <= '1';
SYNTHESIZED_WIRE_116 <= '1';
SYNTHESIZED_WIRE_117 <= '1';



b2v_inst : 74283_0
PORT MAP(CIN => SYNTHESIZED_WIRE_118,
		 A1 => Vaga1,
		 A2 => SYNTHESIZED_WIRE_118,
		 B2 => SYNTHESIZED_WIRE_118,
		 A3 => SYNTHESIZED_WIRE_118,
		 A4 => SYNTHESIZED_WIRE_118,
		 B4 => SYNTHESIZED_WIRE_118,
		 B1 => Vaga2,
		 B3 => SYNTHESIZED_WIRE_118,
		 SUM4 => SYNTHESIZED_WIRE_13,
		 SUM1 => SYNTHESIZED_WIRE_9,
		 SUM2 => SYNTHESIZED_WIRE_10,
		 SUM3 => SYNTHESIZED_WIRE_12);


SYNTHESIZED_WIRE_118 <= NOT(SYNTHESIZED_WIRE_7);







b2v_inst14 : 74283_1
PORT MAP(CIN => SYNTHESIZED_WIRE_118,
		 A1 => SYNTHESIZED_WIRE_9,
		 A2 => SYNTHESIZED_WIRE_10,
		 B2 => SYNTHESIZED_WIRE_118,
		 A3 => SYNTHESIZED_WIRE_12,
		 A4 => SYNTHESIZED_WIRE_13,
		 B4 => SYNTHESIZED_WIRE_118,
		 B1 => Vaga3,
		 B3 => SYNTHESIZED_WIRE_118,
		 SUM4 => SYNTHESIZED_WIRE_21,
		 SUM1 => SYNTHESIZED_WIRE_17,
		 SUM2 => SYNTHESIZED_WIRE_18,
		 SUM3 => SYNTHESIZED_WIRE_20);


b2v_inst15 : 74283_2
PORT MAP(CIN => SYNTHESIZED_WIRE_119,
		 A1 => SYNTHESIZED_WIRE_17,
		 A2 => SYNTHESIZED_WIRE_18,
		 B2 => SYNTHESIZED_WIRE_119,
		 A3 => SYNTHESIZED_WIRE_20,
		 A4 => SYNTHESIZED_WIRE_21,
		 B4 => SYNTHESIZED_WIRE_119,
		 B1 => Vaga4,
		 B3 => SYNTHESIZED_WIRE_119,
		 SUM4 => SYNTHESIZED_WIRE_29,
		 SUM1 => SYNTHESIZED_WIRE_25,
		 SUM2 => SYNTHESIZED_WIRE_26,
		 SUM3 => SYNTHESIZED_WIRE_28);


b2v_inst16 : 74283_3
PORT MAP(CIN => SYNTHESIZED_WIRE_119,
		 A1 => SYNTHESIZED_WIRE_25,
		 A2 => SYNTHESIZED_WIRE_26,
		 B2 => SYNTHESIZED_WIRE_119,
		 A3 => SYNTHESIZED_WIRE_28,
		 A4 => SYNTHESIZED_WIRE_29,
		 B4 => SYNTHESIZED_WIRE_119,
		 B1 => Vaga5,
		 B3 => SYNTHESIZED_WIRE_119,
		 SUM4 => SYNTHESIZED_WIRE_37,
		 SUM1 => SYNTHESIZED_WIRE_33,
		 SUM2 => SYNTHESIZED_WIRE_34,
		 SUM3 => SYNTHESIZED_WIRE_36);


b2v_inst17 : 74283_4
PORT MAP(CIN => SYNTHESIZED_WIRE_120,
		 A1 => SYNTHESIZED_WIRE_33,
		 A2 => SYNTHESIZED_WIRE_34,
		 B2 => SYNTHESIZED_WIRE_120,
		 A3 => SYNTHESIZED_WIRE_36,
		 A4 => SYNTHESIZED_WIRE_37,
		 B4 => SYNTHESIZED_WIRE_120,
		 B1 => Vaga6,
		 B3 => SYNTHESIZED_WIRE_120,
		 SUM4 => SYNTHESIZED_WIRE_45,
		 SUM1 => SYNTHESIZED_WIRE_41,
		 SUM2 => SYNTHESIZED_WIRE_42,
		 SUM3 => SYNTHESIZED_WIRE_44);


b2v_inst18 : 74283_5
PORT MAP(CIN => SYNTHESIZED_WIRE_120,
		 A1 => SYNTHESIZED_WIRE_41,
		 A2 => SYNTHESIZED_WIRE_42,
		 B2 => SYNTHESIZED_WIRE_120,
		 A3 => SYNTHESIZED_WIRE_44,
		 A4 => SYNTHESIZED_WIRE_45,
		 B4 => SYNTHESIZED_WIRE_120,
		 B1 => Vaga7,
		 B3 => SYNTHESIZED_WIRE_120,
		 SUM4 => SYNTHESIZED_WIRE_53,
		 SUM1 => SYNTHESIZED_WIRE_49,
		 SUM2 => SYNTHESIZED_WIRE_50,
		 SUM3 => SYNTHESIZED_WIRE_52);


b2v_inst19 : 74283_6
PORT MAP(CIN => SYNTHESIZED_WIRE_121,
		 A1 => SYNTHESIZED_WIRE_49,
		 A2 => SYNTHESIZED_WIRE_50,
		 B2 => SYNTHESIZED_WIRE_121,
		 A3 => SYNTHESIZED_WIRE_52,
		 A4 => SYNTHESIZED_WIRE_53,
		 B4 => SYNTHESIZED_WIRE_121,
		 B1 => Vaga8,
		 B3 => SYNTHESIZED_WIRE_121,
		 SUM4 => SYNTHESIZED_WIRE_62,
		 SUM1 => SYNTHESIZED_WIRE_58,
		 SUM2 => SYNTHESIZED_WIRE_59,
		 SUM3 => SYNTHESIZED_WIRE_61);


SYNTHESIZED_WIRE_119 <= NOT(SYNTHESIZED_WIRE_56);



b2v_inst20 : 74283_7
PORT MAP(CIN => SYNTHESIZED_WIRE_121,
		 A1 => SYNTHESIZED_WIRE_58,
		 A2 => SYNTHESIZED_WIRE_59,
		 B2 => SYNTHESIZED_WIRE_121,
		 A3 => SYNTHESIZED_WIRE_61,
		 A4 => SYNTHESIZED_WIRE_62,
		 B4 => SYNTHESIZED_WIRE_121,
		 B1 => Vaga9,
		 B3 => SYNTHESIZED_WIRE_121,
		 SUM4 => SYNTHESIZED_WIRE_70,
		 SUM1 => SYNTHESIZED_WIRE_66,
		 SUM2 => SYNTHESIZED_WIRE_67,
		 SUM3 => SYNTHESIZED_WIRE_69);


b2v_inst21 : 74283_8
PORT MAP(CIN => SYNTHESIZED_WIRE_122,
		 A1 => SYNTHESIZED_WIRE_66,
		 A2 => SYNTHESIZED_WIRE_67,
		 B2 => SYNTHESIZED_WIRE_122,
		 A3 => SYNTHESIZED_WIRE_69,
		 A4 => SYNTHESIZED_WIRE_70,
		 B4 => SYNTHESIZED_WIRE_122,
		 B1 => Vaga10,
		 B3 => SYNTHESIZED_WIRE_122,
		 SUM4 => SYNTHESIZED_WIRE_78,
		 SUM1 => SYNTHESIZED_WIRE_74,
		 SUM2 => SYNTHESIZED_WIRE_75,
		 SUM3 => SYNTHESIZED_WIRE_77);


b2v_inst22 : 74283_9
PORT MAP(CIN => SYNTHESIZED_WIRE_122,
		 A1 => SYNTHESIZED_WIRE_74,
		 A2 => SYNTHESIZED_WIRE_75,
		 B2 => SYNTHESIZED_WIRE_122,
		 A3 => SYNTHESIZED_WIRE_77,
		 A4 => SYNTHESIZED_WIRE_78,
		 B4 => SYNTHESIZED_WIRE_122,
		 B1 => Vaga11,
		 B3 => SYNTHESIZED_WIRE_122,
		 SUM4 => SYNTHESIZED_WIRE_86,
		 SUM1 => SYNTHESIZED_WIRE_82,
		 SUM2 => SYNTHESIZED_WIRE_83,
		 SUM3 => SYNTHESIZED_WIRE_85);


b2v_inst23 : 74283_10
PORT MAP(CIN => SYNTHESIZED_WIRE_123,
		 A1 => SYNTHESIZED_WIRE_82,
		 A2 => SYNTHESIZED_WIRE_83,
		 B2 => SYNTHESIZED_WIRE_123,
		 A3 => SYNTHESIZED_WIRE_85,
		 A4 => SYNTHESIZED_WIRE_86,
		 B4 => SYNTHESIZED_WIRE_123,
		 B1 => Vaga12,
		 B3 => SYNTHESIZED_WIRE_123,
		 SUM4 => SYNTHESIZED_WIRE_94,
		 SUM1 => SYNTHESIZED_WIRE_90,
		 SUM2 => SYNTHESIZED_WIRE_91,
		 SUM3 => SYNTHESIZED_WIRE_93);


b2v_inst24 : 74283_11
PORT MAP(CIN => SYNTHESIZED_WIRE_123,
		 A1 => SYNTHESIZED_WIRE_90,
		 A2 => SYNTHESIZED_WIRE_91,
		 B2 => SYNTHESIZED_WIRE_123,
		 A3 => SYNTHESIZED_WIRE_93,
		 A4 => SYNTHESIZED_WIRE_94,
		 B4 => SYNTHESIZED_WIRE_123,
		 B1 => Vaga13,
		 B3 => SYNTHESIZED_WIRE_123,
		 SUM4 => SYNTHESIZED_WIRE_102,
		 SUM1 => SYNTHESIZED_WIRE_98,
		 SUM2 => SYNTHESIZED_WIRE_99,
		 SUM3 => SYNTHESIZED_WIRE_101);


b2v_inst25 : 74283_12
PORT MAP(CIN => SYNTHESIZED_WIRE_124,
		 A1 => SYNTHESIZED_WIRE_98,
		 A2 => SYNTHESIZED_WIRE_99,
		 B2 => SYNTHESIZED_WIRE_124,
		 A3 => SYNTHESIZED_WIRE_101,
		 A4 => SYNTHESIZED_WIRE_102,
		 B4 => SYNTHESIZED_WIRE_124,
		 B1 => Vaga14,
		 B3 => SYNTHESIZED_WIRE_124,
		 SUM4 => SYNTHESIZED_WIRE_110,
		 SUM1 => SYNTHESIZED_WIRE_106,
		 SUM2 => SYNTHESIZED_WIRE_107,
		 SUM3 => SYNTHESIZED_WIRE_109);


b2v_inst26 : 74283_13
PORT MAP(CIN => SYNTHESIZED_WIRE_124,
		 A1 => SYNTHESIZED_WIRE_106,
		 A2 => SYNTHESIZED_WIRE_107,
		 B2 => SYNTHESIZED_WIRE_124,
		 A3 => SYNTHESIZED_WIRE_109,
		 A4 => SYNTHESIZED_WIRE_110,
		 B4 => SYNTHESIZED_WIRE_124,
		 B1 => Vaga15,
		 B3 => SYNTHESIZED_WIRE_124,
		 SUM4 => pin_name4,
		 SUM1 => pin_name1,
		 SUM2 => pin_name2,
		 SUM3 => pin_name3);



SYNTHESIZED_WIRE_120 <= NOT(SYNTHESIZED_WIRE_113);



SYNTHESIZED_WIRE_121 <= NOT(SYNTHESIZED_WIRE_114);



SYNTHESIZED_WIRE_122 <= NOT(SYNTHESIZED_WIRE_115);



SYNTHESIZED_WIRE_123 <= NOT(SYNTHESIZED_WIRE_116);



SYNTHESIZED_WIRE_124 <= NOT(SYNTHESIZED_WIRE_117);





END bdf_type;